`ifndef __CPU_ENDIANESS_VH__
`define __CPU_ENDIANESS_VH__

`define BigEndianCPU 1'b0

`endif
