`define HAS_CACHE
`define PERF_COUNTER
