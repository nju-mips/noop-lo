`define SRAMLIKE_IF
